`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/26/2025 11:25:06 AM
// Design Name: 
// Module Name: Parity_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Parity_tb();
  reg [3:0]b;
  wire p;
  Even_Parity_4bit DUT(b,p);
  
  initial
  begin
   $dumpfile("Even_Parity_4bit.vcd");
   $dumpvars(0,Parity_tb);
   $monitor($time,"b=%b,p=%b",b,p);
   
   #5 b=4'b0000;
   #5 b=4'b0001;
   #5 b=4'b0010;
   #5 b=4'b0011;
   #5 b=4'b0100; 
   #5 b=4'b0101;
   #5 b=4'b0110;
   #5 b=4'b0111;
   #5 b=4'b1000;
   #5 b=4'b1001;
   #5 b=4'b1010;
   #5 b=4'b1011;
   #5 b=4'b1100;
   #5 b=4'b1101;
   #5 b=4'b1110;
   #5 b=4'b1111;
   
   #5 $finish;
    
  end
endmodule
