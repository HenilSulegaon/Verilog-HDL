`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/13/2025 09:34:39 AM
// Design Name: 
// Module Name: binary_2_gray_4bit
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module binary_2_gray_4bit(B,G);
 input [3:0] B;
 output [3:0] G;
 
 assign G[3]=B[3];
 assign G[2]=B[2]^B[3];
 assign G[1]=B[1]^B[2];
 assign G[0]=B[0]^B[1];
endmodule
