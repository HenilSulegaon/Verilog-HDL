`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/16/2025 10:19:15 AM
// Design Name: 
// Module Name: message_print1
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


//module message_print1();
  
//endmodule



module message_print1();
  reg [0:6]a;
  reg [0:6]b;
  reg [0:6]c;
  reg [0:14]r;
  
  initial
  begin
     
     {a[0],a[1],a[2],a[3],a[4],a[5],a[6]} = 7'b1111111; #10;
     {a[0],a[1],a[2],a[3],a[4],a[5],a[6]} = 7'b0001000; #10;
     {a[0],a[1],a[2],a[3],a[4],a[5],a[6]} = 7'b0001000; #10;  // H  
     {a[0],a[1],a[2],a[3],a[4],a[5],a[6]} = 7'b0001000; #10;
     {a[0],a[1],a[2],a[3],a[4],a[5],a[6]} = 7'b1111111; #10;
     
     {a[0],a[1],a[2],a[3],a[4],a[5],a[6]} = 7'b0000000; #10;
     
     {a[0],a[1],a[2],a[3],a[4],a[5],a[6]} = 7'b1111111; #10;
     {a[0],a[1],a[2],a[3],a[4],a[5],a[6]} = 7'b1001001; #10;
     {a[0],a[1],a[2],a[3],a[4],a[5],a[6]} = 7'b1001001; #10; // E
     {a[0],a[1],a[2],a[3],a[4],a[5],a[6]} = 7'b1001001; #10;
     
     {a[0],a[1],a[2],a[3],a[4],a[5],a[6]} = 7'b0000000; #10;
     
     {a[0],a[1],a[2],a[3],a[4],a[5],a[6]} = 7'b1111111; #10;
     {a[0],a[1],a[2],a[3],a[4],a[5],a[6]} = 7'b0000001; #10;
     {a[0],a[1],a[2],a[3],a[4],a[5],a[6]} = 7'b0000001; #10;  // L
     {a[0],a[1],a[2],a[3],a[4],a[5],a[6]} = 7'b0000001; #10;
     
     {a[0],a[1],a[2],a[3],a[4],a[5],a[6]} = 7'b0000000; #10;
     
     {a[0],a[1],a[2],a[3],a[4],a[5],a[6]} = 7'b1111111; #10;
     {a[0],a[1],a[2],a[3],a[4],a[5],a[6]} = 7'b0000001; #10;
     {a[0],a[1],a[2],a[3],a[4],a[5],a[6]} = 7'b0000001; #10;  // L
     {a[0],a[1],a[2],a[3],a[4],a[5],a[6]} = 7'b0000001; #10;
     
     
     {a[0],a[1],a[2],a[3],a[4],a[5],a[6]} = 7'b0000000; #10;
     
     {a[0],a[1],a[2],a[3],a[4],a[5],a[6]} = 7'b1111111; #10;
     {a[0],a[1],a[2],a[3],a[4],a[5],a[6]} = 7'b1000001; #10;
     {a[0],a[1],a[2],a[3],a[4],a[5],a[6]} = 7'b1000001; #10;  // O
     {a[0],a[1],a[2],a[3],a[4],a[5],a[6]} = 7'b1000001; #10;
     {a[0],a[1],a[2],a[3],a[4],a[5],a[6]} = 7'b1111111; #10;
     
     {a[0],a[1],a[2],a[3],a[4],a[5],a[6]} = 7'b0000000; #10;
//     $finish;
  end
  
  initial
  begin
     {b[0],b[1],b[2],b[3],b[4],b[5],b[6]} = 7'b1111111; #10;
     {b[0],b[1],b[2],b[3],b[4],b[5],b[6]} = 7'b1000001; #10;
     {b[0],b[1],b[2],b[3],b[4],b[5],b[6]} = 7'b1000001; #10;
     {b[0],b[1],b[2],b[3],b[4],b[5],b[6]} = 7'b1000101; #10; // G
     {b[0],b[1],b[2],b[3],b[4],b[5],b[6]} = 7'b1000101; #10;
     {b[0],b[1],b[2],b[3],b[4],b[5],b[6]} = 7'b1000111; #10;
     
     {b[0],b[1],b[2],b[3],b[4],b[5],b[6]} = 7'b0000000; #10;
     
     {b[0],b[1],b[2],b[3],b[4],b[5],b[6]} = 7'b1111111; #10;
     {b[0],b[1],b[2],b[3],b[4],b[5],b[6]} = 7'b1000001; #10;
     {b[0],b[1],b[2],b[3],b[4],b[5],b[6]} = 7'b1000001; #10;
     {b[0],b[1],b[2],b[3],b[4],b[5],b[6]} = 7'b1000001; #10; // O
     {b[0],b[1],b[2],b[3],b[4],b[5],b[6]} = 7'b1111111; #10;
     
     {b[0],b[1],b[2],b[3],b[4],b[5],b[6]} = 7'b0000000; #10;
     
     {b[0],b[1],b[2],b[3],b[4],b[5],b[6]} = 7'b1111111; #10;
     {b[0],b[1],b[2],b[3],b[4],b[5],b[6]} = 7'b1000001; #10;
     {b[0],b[1],b[2],b[3],b[4],b[5],b[6]} = 7'b1000001; #10;
     {b[0],b[1],b[2],b[3],b[4],b[5],b[6]} = 7'b1000001; #10; // O
     {b[0],b[1],b[2],b[3],b[4],b[5],b[6]} = 7'b1111111; #10;
     
     {b[0],b[1],b[2],b[3],b[4],b[5],b[6]} = 7'b0000000; #10;
     
     {b[0],b[1],b[2],b[3],b[4],b[5],b[6]} = 7'b1111111; #10;
     {b[0],b[1],b[2],b[3],b[4],b[5],b[6]} = 7'b1000001; #10;
     {b[0],b[1],b[2],b[3],b[4],b[5],b[6]} = 7'b0100010; #10;  // D
     {b[0],b[1],b[2],b[3],b[4],b[5],b[6]} = 7'b0011100; #10;
     
     {b[0],b[1],b[2],b[3],b[4],b[5],b[6]} = 7'b0000000; #10;
//     $finish;
  end
  
  initial
  begin
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b1111111; #10;
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b0100000; #10;
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b0010000; #10;
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b0001000; #10;  // M
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b0010000; #10;
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b0100000; #10;
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b1111111; #10;
    
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b0000000; #10;
    
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b1111111; #10;
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b1000001; #10;
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b1000001; #10;  // O
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b1000001; #10;
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b1111111; #10;
    
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b0000000; #10;
    
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b1111111; #10;
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b1001100; #10;
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b1001010; #10;  // R
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b1001001; #10;
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b1111001; #10;
    
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b0000000; #10;
    
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b1111111; #10;
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b0100000; #10;
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b0010000; #10;
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b0001000; #10;  // N
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b0000100; #10;
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b0000010; #10;
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b1111111; #10;
    
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b0000000; #10;
    
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b1000001; #10;
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b1000001; #10;
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b1111111; #10;  // I
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b1000001; #10;
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b1000001; #10;
    
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b0000000; #10;
    
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b1111111; #10;
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b0100000; #10;
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b0010000; #10;
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b0001000; #10;  // N
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b0000100; #10;
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b0000010; #10;
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b1111111; #10;
    
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b0000000; #10;
    
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b1111111; #10;
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b1000001; #10;
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b1000001; #10;
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b1000101; #10;  // G
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b1000101; #10;
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b1000111; #10;
    
    {c[0],c[1],c[2],c[3],c[4],c[5],c[6]}= 7'b0000000; #10;
//    $finish;
  end
  
  initial
  begin
    
    {r[0], r[1], r[2], r[3], r[4], r[5], r[6],r[7],r[8],r[9],r[10],r[11],r[12],r[13],r[14]} =15'b000000000000000; #20;
    {r[0], r[1], r[2], r[3], r[4], r[5], r[6],r[7],r[8],r[9],r[10],r[11],r[12],r[13],r[14]} =15'b000000000000000; #20;
    {r[0], r[1], r[2], r[3], r[4], r[5], r[6],r[7],r[8],r[9],r[10],r[11],r[12],r[13],r[14]} =15'b000000000000000; #20;
    {r[0], r[1], r[2], r[3], r[4], r[5], r[6],r[7],r[8],r[9],r[10],r[11],r[12],r[13],r[14]} =15'b000000000000000; #20;
    {r[0], r[1], r[2], r[3], r[4], r[5], r[6],r[7],r[8],r[9],r[10],r[11],r[12],r[13],r[14]} =15'b000000000000000; #20;
    
    {r[0], r[1], r[2], r[3], r[4], r[5], r[6],r[7],r[8],r[9],r[10],r[11],r[12],r[13],r[14]} = 15'b111111111111111; #5;  //c1
    {r[0], r[1], r[2], r[3], r[4], r[5], r[6],r[7],r[8],r[9],r[10],r[11],r[12],r[13],r[14]} = 15'b100000000000001; #5;  // c2
    {r[0], r[1], r[2], r[3], r[4], r[5], r[6],r[7],r[8],r[9],r[10],r[11],r[12],r[13],r[14]} = 15'b100010000000001; #5;  //c3
    {r[0], r[1], r[2], r[3], r[4], r[5], r[6],r[7],r[8],r[9],r[10],r[11],r[12],r[13],r[14]} = 15'b100101000000001; #5;
    {r[0], r[1], r[2], r[3], r[4], r[5], r[6],r[7],r[8],r[9],r[10],r[11],r[12],r[13],r[14]} = 15'b101000100000001; #5;
    {r[0], r[1], r[2], r[3], r[4], r[5], r[6],r[7],r[8],r[9],r[10],r[11],r[12],r[13],r[14]} = 15'b100101000000001; #5;
    {r[0], r[1], r[2], r[3], r[4], r[5], r[6],r[7],r[8],r[9],r[10],r[11],r[12],r[13],r[14]} = 15'b100010000000001; #5;
    {r[0], r[1], r[2], r[3], r[4], r[5], r[6],r[7],r[8],r[9],r[10],r[11],r[12],r[13],r[14]} = 15'b100000000110001; #5;
    {r[0], r[1], r[2], r[3], r[4], r[5], r[6],r[7],r[8],r[9],r[10],r[11],r[12],r[13],r[14]} = 15'b100000000101001; #5;
    {r[0], r[1], r[2], r[3], r[4], r[5], r[6],r[7],r[8],r[9],r[10],r[11],r[12],r[13],r[14]} = 15'b100000000100101; #5;
    {r[0], r[1], r[2], r[3], r[4], r[5], r[6],r[7],r[8],r[9],r[10],r[11],r[12],r[13],r[14]} = 15'b100000000101001; #5;
    {r[0], r[1], r[2], r[3], r[4], r[5], r[6],r[7],r[8],r[9],r[10],r[11],r[12],r[13],r[14]} = 15'b100000000110001; #5;  // Smile 
    {r[0], r[1], r[2], r[3], r[4], r[5], r[6],r[7],r[8],r[9],r[10],r[11],r[12],r[13],r[14]} = 15'b100010000000001; #5;
    {r[0], r[1], r[2], r[3], r[4], r[5], r[6],r[7],r[8],r[9],r[10],r[11],r[12],r[13],r[14]} = 15'b100101000000001; #5;
    {r[0], r[1], r[2], r[3], r[4], r[5], r[6],r[7],r[8],r[9],r[10],r[11],r[12],r[13],r[14]} = 15'b101000100000001; #5;
    {r[0], r[1], r[2], r[3], r[4], r[5], r[6],r[7],r[8],r[9],r[10],r[11],r[12],r[13],r[14]} = 15'b100101000000001; #5;
    {r[0], r[1], r[2], r[3], r[4], r[5], r[6],r[7],r[8],r[9],r[10],r[11],r[12],r[13],r[14]} = 15'b100010000000001; #5;
    {r[0], r[1], r[2], r[3], r[4], r[5], r[6],r[7],r[8],r[9],r[10],r[11],r[12],r[13],r[14]} = 15'b100000000000001; #5;
    {r[0], r[1], r[2], r[3], r[4], r[5], r[6],r[7],r[8],r[9],r[10],r[11],r[12],r[13],r[14]} = 15'b111111111111111; #5;
    
     {r[0], r[1], r[2], r[3], r[4], r[5], r[6],r[7],r[8],r[9],r[10],r[11],r[12],r[13],r[14]} =15'b000000000000000; #5;
//    $finish;
  end
endmodule