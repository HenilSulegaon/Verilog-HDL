`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/13/2025 09:38:41 AM
// Design Name: 
// Module Name: binary_2_gray_4bit_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module binary_2_gray_4bit_tb();
  reg [3:0]B;
  wire [3:0]G;
  binary_2_gray_4bit DUT(B,G);
  
  initial
  begin
    $dumpfile("binary_2_gray_4bit.vcd");
    $dumpvars(0,binary_2_gray_4bit_tb);
    $monitor($time,"B=%b,G=%b",B,G);
    
    #5 B=4'b0000;
    #5 B=4'b0001;
    #5 B=4'b0010;
    #5 B=4'b0011;
    #5 B=4'b0100;
    #5 B=4'b0101;
    #5 B=4'b0110;
    #5 B=4'b0111;
    #5 B=4'b1000;
    #5 B=4'b1001;
    #5 B=4'b1010;
    #5 B=4'b1011;
    #5 B=4'b1100;
    #5 B=4'b1101;
    #5 B=4'b1110;
    #5 B=4'b1111;
    #5 $finish;
    
  end
endmodule
